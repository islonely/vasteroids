module main

import gg
import net

fn (mut app App) draw_multiplayer_in_game() {
}

fn (mut app App) update_multiplayer_in_game() {
}
